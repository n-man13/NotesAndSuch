module Adder_4_tb;
    reg [3:0] a;
    reg [3:0] b;
    reg [4:0] s;
    integer i;

    FourBitAdder four(a, b, s);

    initial begin
        a = 4'b0000;
        b = 4'b0000;
        for (i = 0; i < 16; i = i + 1) begin
            a = i;
            for (integer j = 0; j < 16; j = j + 1) begin
                b = j;
            end
            #10
        end
    end

    initial begin
        $dumpfile("test_four.vcd");
        $dumpvars(0,Adder_4_tb);
    end

endmodule